module main

fn main() {
	println([9,8,7,6,5,4,3,2,1].sorted())
}